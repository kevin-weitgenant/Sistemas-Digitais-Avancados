library verilog;
use verilog.vl_types.all;
entity mux8pra1_vlg_vec_tst is
end mux8pra1_vlg_vec_tst;
