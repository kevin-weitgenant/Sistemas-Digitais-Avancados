library verilog;
use verilog.vl_types.all;
entity mux2pra1_vlg_vec_tst is
end mux2pra1_vlg_vec_tst;
