library verilog;
use verilog.vl_types.all;
entity ULA1_vlg_vec_tst is
end ULA1_vlg_vec_tst;
