library verilog;
use verilog.vl_types.all;
entity ULA2_vlg_vec_tst is
end ULA2_vlg_vec_tst;
