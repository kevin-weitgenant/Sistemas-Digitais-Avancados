library verilog;
use verilog.vl_types.all;
entity somador_subtrator_nbits_vlg_vec_tst is
end somador_subtrator_nbits_vlg_vec_tst;
